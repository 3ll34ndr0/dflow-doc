magic
tech scmos
magscale 1 2
timestamp 1429114932
<< checkpaint >>
rect -78 -66 150 270
<< nwell >>
rect -18 96 90 210
<< ntransistor >>
rect 14 12 18 52
rect 30 12 34 52
rect 46 12 50 52
rect 62 12 66 52
<< ptransistor >>
rect 14 108 18 188
rect 30 108 34 188
rect 46 108 50 188
rect 62 108 66 188
<< ndiffusion >>
rect 4 51 14 52
rect 12 13 14 51
rect 4 12 14 13
rect 18 51 30 52
rect 18 13 20 51
rect 28 13 30 51
rect 18 12 30 13
rect 34 51 46 52
rect 34 13 36 51
rect 44 13 46 51
rect 34 12 46 13
rect 50 51 62 52
rect 50 13 52 51
rect 60 13 62 51
rect 50 12 62 13
rect 66 51 76 52
rect 66 13 68 51
rect 66 12 76 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 109 14 187
rect 4 108 14 109
rect 18 187 30 188
rect 18 109 20 187
rect 28 109 30 187
rect 18 108 30 109
rect 34 187 46 188
rect 34 109 36 187
rect 44 109 46 187
rect 34 108 46 109
rect 50 187 62 188
rect 50 109 52 187
rect 60 109 62 187
rect 50 108 62 109
rect 66 187 76 188
rect 66 109 68 187
rect 66 108 76 109
<< ndcontact >>
rect 4 13 12 51
rect 20 13 28 51
rect 36 13 44 51
rect 52 13 60 51
rect 68 13 76 51
<< pdcontact >>
rect 4 109 12 187
rect 20 109 28 187
rect 36 109 44 187
rect 52 109 60 187
rect 68 109 76 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
rect 60 -4 68 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
rect 60 196 68 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 46 188 50 192
rect 62 188 66 192
rect 14 106 18 108
rect 30 106 34 108
rect 46 106 50 108
rect 62 106 66 108
rect 14 102 66 106
rect 14 66 18 102
rect 12 60 18 66
rect 12 58 66 60
rect 14 56 66 58
rect 14 52 18 56
rect 30 52 34 56
rect 46 52 50 56
rect 62 52 66 56
rect 14 8 18 12
rect 30 8 34 12
rect 46 8 50 12
rect 62 8 66 12
<< polycontact >>
rect 4 58 12 66
<< metal1 >>
rect -4 204 84 206
rect 4 196 28 204
rect 36 196 60 204
rect 68 196 84 204
rect -4 194 84 196
rect 4 187 12 194
rect 4 108 12 109
rect 20 187 28 188
rect 20 102 28 109
rect 36 187 44 194
rect 36 108 44 109
rect 52 187 60 188
rect 52 102 60 109
rect 68 187 76 194
rect 68 108 76 109
rect 20 94 60 102
rect 4 66 12 74
rect 52 66 60 94
rect 20 58 60 66
rect 4 51 12 52
rect 4 6 12 13
rect 20 51 28 58
rect 20 12 28 13
rect 36 51 44 52
rect 36 6 44 13
rect 52 51 60 58
rect 52 12 60 13
rect 68 51 76 52
rect 68 6 76 13
rect -4 4 84 6
rect 4 -4 28 4
rect 36 -4 60 4
rect 68 -4 84 4
rect -4 -6 84 -4
<< m1p >>
rect 52 86 60 94
rect 4 66 12 74
<< labels >>
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 70 8 70 4 A
rlabel metal1 56 90 56 90 4 Y
<< end >>
