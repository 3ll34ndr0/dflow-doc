magic
tech scmos
magscale 1 2
timestamp 1429114932
<< checkpaint >>
rect -74 -66 138 270
<< nwell >>
rect -14 96 78 210
<< ntransistor >>
rect 20 12 24 52
rect 30 12 34 52
rect 46 12 50 32
<< ptransistor >>
rect 14 108 18 188
rect 30 108 34 188
rect 46 108 50 188
<< ndiffusion >>
rect 10 51 20 52
rect 18 13 20 51
rect 10 12 20 13
rect 24 12 30 52
rect 34 51 44 52
rect 34 13 36 51
rect 44 13 46 32
rect 34 12 46 13
rect 50 31 60 32
rect 50 13 52 31
rect 50 12 60 13
<< pdiffusion >>
rect 4 185 14 188
rect 12 117 14 185
rect 4 108 14 117
rect 18 120 20 188
rect 28 120 30 188
rect 18 108 30 120
rect 34 187 46 188
rect 34 109 36 187
rect 44 109 46 187
rect 34 108 46 109
rect 50 187 60 188
rect 50 109 52 187
rect 50 108 60 109
<< ndcontact >>
rect 10 13 18 51
rect 36 13 44 51
rect 52 13 60 31
<< pdcontact >>
rect 4 117 12 185
rect 20 120 28 188
rect 36 109 44 187
rect 52 109 60 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 46 188 50 192
rect 14 98 18 108
rect 8 58 12 94
rect 30 82 34 108
rect 28 74 34 82
rect 8 54 24 58
rect 20 52 24 54
rect 30 52 34 74
rect 46 32 50 108
rect 20 8 24 12
rect 30 8 34 12
rect 46 8 50 12
<< polycontact >>
rect 12 90 20 98
rect 20 74 28 82
rect 50 38 58 46
<< metal1 >>
rect -4 204 68 206
rect 4 196 28 204
rect 36 196 68 204
rect -4 194 68 196
rect 20 188 28 194
rect 4 185 12 188
rect 36 187 44 188
rect 4 114 12 117
rect 4 109 36 114
rect 4 108 44 109
rect 52 187 60 188
rect 52 108 60 109
rect 4 90 12 94
rect 52 94 58 108
rect 4 88 20 90
rect 36 88 60 94
rect 4 86 12 88
rect 20 66 28 74
rect 36 52 42 88
rect 52 86 60 88
rect 10 51 18 52
rect 10 6 18 13
rect 36 51 44 52
rect 52 46 60 54
rect 36 12 44 13
rect 52 31 60 32
rect 52 6 60 13
rect -4 4 68 6
rect 4 -4 28 4
rect 36 -4 68 4
rect -4 -6 68 -4
<< m1p >>
rect 4 86 12 94
rect 52 86 60 94
rect 20 66 28 74
rect 52 46 60 54
<< labels >>
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 90 8 90 4 A
rlabel metal1 24 70 24 70 4 B
rlabel metal1 56 90 56 90 4 Y
rlabel metal1 56 50 56 50 4 C
<< end >>
