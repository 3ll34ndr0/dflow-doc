magic
tech scmos
magscale 1 2
timestamp 1429114932
<< checkpaint >>
rect -76 -66 152 270
<< nwell >>
rect -16 96 92 210
<< ntransistor >>
rect 18 12 22 52
rect 28 12 32 52
rect 52 12 56 52
rect 62 12 66 52
<< ptransistor >>
rect 14 108 18 188
rect 30 108 34 188
rect 46 108 50 188
rect 62 108 66 188
<< ndiffusion >>
rect 8 51 18 52
rect 16 13 18 51
rect 8 12 18 13
rect 22 12 28 52
rect 32 51 52 52
rect 32 13 38 51
rect 46 13 52 51
rect 32 12 52 13
rect 56 12 62 52
rect 66 51 76 52
rect 66 13 68 51
rect 66 12 76 13
<< pdiffusion >>
rect 4 185 14 188
rect 12 117 14 185
rect 4 108 14 117
rect 18 120 20 188
rect 28 120 30 188
rect 18 108 30 120
rect 34 187 46 188
rect 34 109 36 187
rect 44 109 46 187
rect 34 108 46 109
rect 50 176 62 188
rect 50 108 52 176
rect 60 108 62 176
rect 66 187 76 188
rect 66 109 68 187
rect 66 108 76 109
<< ndcontact >>
rect 8 13 16 51
rect 38 13 46 51
rect 68 13 76 51
<< pdcontact >>
rect 4 117 12 185
rect 20 120 28 188
rect 36 109 44 187
rect 52 108 60 176
rect 68 109 76 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
rect 60 -4 68 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
rect 60 196 68 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 46 188 50 192
rect 62 188 66 192
rect 14 98 18 108
rect 30 106 34 108
rect 28 102 34 106
rect 8 58 12 94
rect 8 54 22 58
rect 18 52 22 54
rect 28 52 32 102
rect 46 80 50 108
rect 62 106 66 108
rect 62 102 70 106
rect 66 94 68 102
rect 48 78 50 80
rect 48 58 52 78
rect 66 62 70 94
rect 62 58 70 62
rect 48 54 56 58
rect 52 52 56 54
rect 62 52 66 58
rect 18 8 22 12
rect 28 8 32 12
rect 52 8 56 12
rect 62 8 66 12
<< polycontact >>
rect 12 90 20 98
rect 20 74 28 82
rect 68 94 76 102
rect 50 78 58 86
<< metal1 >>
rect -4 204 84 206
rect 4 196 28 204
rect 36 196 60 204
rect 68 196 84 204
rect -4 194 84 196
rect 20 188 28 194
rect 4 185 12 188
rect 36 187 76 188
rect 4 114 12 117
rect 4 109 36 114
rect 44 182 68 187
rect 4 108 44 109
rect 68 108 76 109
rect 52 102 58 108
rect 4 90 12 94
rect 38 96 58 102
rect 38 94 44 96
rect 4 88 20 90
rect 4 86 12 88
rect 36 86 44 94
rect 68 86 76 94
rect 20 66 28 74
rect 38 52 44 86
rect 52 74 58 78
rect 52 66 60 74
rect 8 51 16 52
rect 8 6 16 13
rect 34 51 50 52
rect 34 13 38 51
rect 46 13 50 51
rect 34 12 50 13
rect 68 51 76 52
rect 68 6 76 13
rect -4 4 84 6
rect 4 -4 28 4
rect 36 -4 60 4
rect 68 -4 84 4
rect -4 -6 84 -4
<< m1p >>
rect 4 86 12 94
rect 36 86 44 94
rect 68 86 76 94
rect 20 66 28 74
rect 52 66 60 74
<< labels >>
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 72 90 72 90 4 C
rlabel metal1 56 70 56 70 4 D
rlabel metal1 40 90 40 90 4 Y
rlabel metal1 8 90 8 90 4 A
rlabel metal1 24 70 24 70 4 B
<< end >>
